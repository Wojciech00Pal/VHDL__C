library IEEE; 
use IEEE.STD_LOGIC_1164.ALL;

entity serializer_tb is 
end serializer_tb;


architecture TEST of serializer_tb is